module prng(
    input clk, // Входной сигнал тактового генератора
//    input rst, // Входной сигнал сброса
    output reg [7:0] out // Выходной 8-битный регистр
);

// Внутренний 8-битный регистр для хранения текущего состояния
reg [7:0] state;

// При каждом такте обновляем состояние и выход по формуле x[n+1] = (a * x[n] + c) mod m
always @(posedge clk) begin
    state <= (8'b00011101 ^ state ^ 8'b01110001) % 9'b100000000;
    out <= state;
end

endmodule