//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.9 Beta-6
//Part Number: GW1NSR-LV4CQN48PC7/I6
//Device: GW1NSR-4C
//Created Time: Tue Nov 14 23:51:50 2023

module Gowin_pROM (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [10:0] ad;

wire [23:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 8;
defparam prom_inst_0.RESET_MODE = "ASYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h8C31E1B9095DE0A02FF1F4E39F88A69CB04DF99223AAEB52606FAB92FECD6BFF;
defparam prom_inst_0.INIT_RAM_01 = 256'h2AE19E9DA6974851094176CA0A771CDB3A277C953FE005689ACE47992BD4DF65;
defparam prom_inst_0.INIT_RAM_02 = 256'h4A736A032BE34AD4429288D6B771F5A3A35ACBD1184131AEC922DD632DB73614;
defparam prom_inst_0.INIT_RAM_03 = 256'h5D4E049113930AA12703F796CB03D2CC6AC886E2EADBDC1936C2E30394195992;
defparam prom_inst_0.INIT_RAM_04 = 256'h1150C0244F433D2C5E88C2533337881F7FB8EFD9EC2CF657DBDD64311AB03FE8;
defparam prom_inst_0.INIT_RAM_05 = 256'h7B5655E98C32952C038BEE0EB2F153606F8179030E71CE5829966CDBC899C368;
defparam prom_inst_0.INIT_RAM_06 = 256'hC8C085A6A0525BBB59CF8B2EAC336172D8F5721CFCC1A251669F382E3FCF0292;
defparam prom_inst_0.INIT_RAM_07 = 256'h742907B797DD3567A684623F0A9D5FA91599B7A6EE8B96D91108CCC11BE9A467;
defparam prom_inst_0.INIT_RAM_08 = 256'hA2807F061267AAB38ED526DC3634496DBD2BCD039A2517A996B68EB078DBECC6;
defparam prom_inst_0.INIT_RAM_09 = 256'h0A5E8669200CC98C49F51561600F3B2F6FE470F4B3872133339DEF0BCCC10245;
defparam prom_inst_0.INIT_RAM_0A = 256'h4B048D27031F77E573351744766DC000CD22B923BA80C2BAA518DA607247B256;
defparam prom_inst_0.INIT_RAM_0B = 256'hAA7056384540C59613878C8D2F39CDD46799EF19E88E634522C9A74C1A32A781;
defparam prom_inst_0.INIT_RAM_0C = 256'h58CBF9DA190B8B7F4DCD4547FD9446AC5F72F2DC3A44B11C3EB28221C5992155;
defparam prom_inst_0.INIT_RAM_0D = 256'h03B163E2880722D47F0219C18BE4F0AD478F5DDE3A93081F1B953C0914625E4B;
defparam prom_inst_0.INIT_RAM_0E = 256'hDB7DC6C407072E0788CF8009ADF1340A6028941D0A0BA5ECBE2CDF7EAEFBE73D;
defparam prom_inst_0.INIT_RAM_0F = 256'h8E848F87EB6DA573CBE11A1C5C368D01D22429CBED9DAB511EF94AA4C93BB566;
defparam prom_inst_0.INIT_RAM_10 = 256'h3760A3A329006182EF76DBBC6180129E2E8A31DD2CBFC91BA6DC81D5F1AEDE79;
defparam prom_inst_0.INIT_RAM_11 = 256'h445ABAB4DBAF829A6DE7DC479B40F9ED4AAA20DBAC960F5458133DD628173B08;
defparam prom_inst_0.INIT_RAM_12 = 256'h45816DE1C8C96875AC5D4F79F35370AC9A68EE7D6C2FBD67D76ED47822056197;
defparam prom_inst_0.INIT_RAM_13 = 256'h06713DA1C07A9C4C633D34CA9F0BE184B2958905359CD346E11BABEBE8A29CC7;
defparam prom_inst_0.INIT_RAM_14 = 256'hF8976B2993DEC2D2ABACA42F2E823CBA6554B1B774B898C4CF4DFC0CF1EE97F2;
defparam prom_inst_0.INIT_RAM_15 = 256'hADD0D7ADA31231E9220393BF5501525FA8876E0F6DFE2BF9E3B4597948C07C24;
defparam prom_inst_0.INIT_RAM_16 = 256'h35A9603CFDDEB3568A3EDE2B39DC157A6F0B814855D690E7AE208A9003551536;
defparam prom_inst_0.INIT_RAM_17 = 256'h082981A2A1AFEAC11CDAE7155FC9AF683F2838433C6D063C23CBDD7DB074D697;
defparam prom_inst_0.INIT_RAM_18 = 256'h7DCADB89C4B7124220B4E4062041E86D194AD94E9130C7BAEDF74DE3E021A8BB;
defparam prom_inst_0.INIT_RAM_19 = 256'hB65473AA04B806016419139C6EBF1644CFB3DB51A6AF2A9B03789A52544E36EA;
defparam prom_inst_0.INIT_RAM_1A = 256'h0EF6616EC99D5B8728167D4D1B002A569D6708DF8124AC3BF3A13D8F83EBFC15;
defparam prom_inst_0.INIT_RAM_1B = 256'h630B83B3577128E90A6B9E9C5BAE108BBE272FF5D5B82E6B472207832C3F0187;
defparam prom_inst_0.INIT_RAM_1C = 256'hF5CCB1A7E1C00149C8C275592A848A2F5AB8806DA51D9E5E05F3FE61B67350F2;
defparam prom_inst_0.INIT_RAM_1D = 256'hCAC4140D95D4A2B3ABE8289D1240D0C4B4D6D3EDE4BE9BE545437E0BBDB6FDCE;
defparam prom_inst_0.INIT_RAM_1E = 256'h2641D706B1D8D33A364B13A0D377DCBF7A222D9E659B88B6B3C760DF1F6D6D1D;
defparam prom_inst_0.INIT_RAM_1F = 256'h9A82C6FBAB372F0181372BC21EF5B37302BB6AB5BEC39D6B9205671C43FB8928;
defparam prom_inst_0.INIT_RAM_20 = 256'h37C338B13BBF48DA22B2765D6546F468848637249E1505A0D2606B9518994947;
defparam prom_inst_0.INIT_RAM_21 = 256'h43ACAFA00039E71FBC547BEFC551E8EC62866E2E49BA65E7EE6E1B5887D2479D;
defparam prom_inst_0.INIT_RAM_22 = 256'hAA78F7E9399CCE14C6E624BBE12D3F41585440AB28A90CE7319D28BAAD0AB6B2;
defparam prom_inst_0.INIT_RAM_23 = 256'hCD3F22EE05AC688F4F8E96CE018E5470900638D9B995B6F3C79BD4CB288FCC21;
defparam prom_inst_0.INIT_RAM_24 = 256'hF308589C5E30ACB21CC9D3622A600AA678F12AC17EE98F888724EF289EF8C9CE;
defparam prom_inst_0.INIT_RAM_25 = 256'h583C43B048D9E0021D1AE5EB990162EB7DD4495AA810781BE8DABE8A14C4745F;
defparam prom_inst_0.INIT_RAM_26 = 256'h014FEFE8D09E5F2326B9E00BBECE7A60DCE799A3AA2F61932F52485370DB7568;
defparam prom_inst_0.INIT_RAM_27 = 256'h32614D347B7662F8ABCE23ED4D84D52C8105BE4541D3DE9C1BADB3B5E710BA36;
defparam prom_inst_0.INIT_RAM_28 = 256'hD80EFE5714EE3942F912E2ACFD2414DEB06D2F5F486DE0BB4E634FD200CA428B;
defparam prom_inst_0.INIT_RAM_29 = 256'hD13FE4C1763EEC27BCD62237C11F14E74B432EC3BE31E2C3D407ABCD41D610B2;
defparam prom_inst_0.INIT_RAM_2A = 256'h0EBC217C3E7BCBAE823DE261B96273B30812C36584B128D3FA91FA3558A28CDF;
defparam prom_inst_0.INIT_RAM_2B = 256'h63B2F81665598631E5D4977013EC2F026EC18903D5FC5D7A43BD190CADB9A4DB;
defparam prom_inst_0.INIT_RAM_2C = 256'hA10E27935C91F01F9551E3E720DCCA1CF46350199A44940E2BAE4BA2F80637FF;
defparam prom_inst_0.INIT_RAM_2D = 256'h724F5BC9B627E5AB27966C5832DD3320FA176105DA7A4BD6CB6BAC0CD6CE13DE;
defparam prom_inst_0.INIT_RAM_2E = 256'hC06FE27BD8193235A162E06FCD0B8A1B3FAA64C2857789790925C9D5D013288B;
defparam prom_inst_0.INIT_RAM_2F = 256'h5CC322239AD5875FAE5DDCC14CD9A863ED0B05648CAD1E2861E17CC86E3D4607;
defparam prom_inst_0.INIT_RAM_30 = 256'hC1646B15D25E1FC192B4012BCA966147272290F498B9EE5A5C6E1AF7F253AB6F;
defparam prom_inst_0.INIT_RAM_31 = 256'hBEBACF4CADDA989C0A2D2564F84DFE664A59744E53ADC42D411F3B04419D09B1;
defparam prom_inst_0.INIT_RAM_32 = 256'h254B388BA3FF7F98F65339E6E90EBF613C7B627432D40A9EE99CD3D46B5A8121;
defparam prom_inst_0.INIT_RAM_33 = 256'h1F826DF8D2832BA9B855EDE25757A72C9423C2EC4731AAEB3CCBBE2F18F936EF;
defparam prom_inst_0.INIT_RAM_34 = 256'hFD93B0AADE891665866B369C154D4367F0E0DC56E100EF3C13A338D01EBBDCB8;
defparam prom_inst_0.INIT_RAM_35 = 256'h53495003B74F04B96FA7EC3270A30C225E88AF9C0E4E7B3DF2FBA96508EE0566;
defparam prom_inst_0.INIT_RAM_36 = 256'hE13202AC92F977FD05109128053BED0F1AA5BECDBD79DBCBB8EA691EA9802CD9;
defparam prom_inst_0.INIT_RAM_37 = 256'h897C3219BE1C2518087D7525221D09F8ED05D0FC7D69120989807B268EFBE618;
defparam prom_inst_0.INIT_RAM_38 = 256'hC7A8C01E29BBBD79A8464D4F875D23A9941EB92E0D278705012C1D77C0A5D2F0;
defparam prom_inst_0.INIT_RAM_39 = 256'hFEAE51AC7FDCC38B05A3D58A9566394ECC6D3025BB9DF744F24B45BAD033E2B6;
defparam prom_inst_0.INIT_RAM_3A = 256'h27CF22F4F8915006828D5333701A810FE2AD002D97517AEF5A9383835EA850B9;
defparam prom_inst_0.INIT_RAM_3B = 256'h2929662EDDE969F1080A5E83FDA21D8DBACBBA49AD1B2222C3E21FC09C0D9536;
defparam prom_inst_0.INIT_RAM_3C = 256'h6C347E8C9E4002FB72BC3305E108A37A574426AE479D30D92B856AAF94D66FFE;
defparam prom_inst_0.INIT_RAM_3D = 256'hC1B76048CFAFD9C10DBFA1B347AF44C52E590C2FAA716DB51D3BF818B71F209D;
defparam prom_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000016AA9AAC886E80AE35621D2DC35265AC;

endmodule //Gowin_pROM
